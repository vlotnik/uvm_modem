`timescale 100ps/100ps

module tb_top;
//--------------------------------------------------------------------------------------------------------------------------------
// libraries
//--------------------------------------------------------------------------------------------------------------------------------
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "common_macros.svh"

    import pkg_modem::*;

    `print_logo

//--------------------------------------------------------------------------------------------------------------------------------
// clock generator
//--------------------------------------------------------------------------------------------------------------------------------
    bit clk = 0;
    // 100 MHz
    always #50 clk = ~clk;

//--------------------------------------------------------------------------------------------------------------------------------
// interface
//--------------------------------------------------------------------------------------------------------------------------------
    if_ddc_bfm #(.INCH_NUMBER(2)) if_ddc_bfm_h();

    assign if_ddc_bfm_h.clk         = clk;
    assign if_ddc_bfm_h.iq_v        = 1;

endmodule