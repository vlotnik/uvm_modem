//--------------------------------------------------------------------------------------------------------------------------------
// name : iqmap
//--------------------------------------------------------------------------------------------------------------------------------
class iqmap extends iqmap_base;
    `uvm_object_utils(iqmap)
    `uvm_object_new

    extern function void init_plane(t_modulation mod);
endclass

//-------------------------------------------------------------------------------------------------------------------------------
// IMPLEMENTATION
//-------------------------------------------------------------------------------------------------------------------------------
function void iqmap::init_plane(t_modulation mod);
    case(mod)
        BPSK : super.plane = {
             0.7070,  0.7070,       // 0
            -0.7070, -0.7070        // 1
        };

        QPSK : super.plane = {
             0.7070,  0.7070,       // 0
             0.7070, -0.7070,       // 1
            -0.7070,  0.7070,       // 2
            -0.7070, -0.7070        // 3
        };

        PSK8 : super.plane = {
             1.0000,  0.0000,       // 0
             0.7070,  0.7070,       // 1
             0.0000,  1.0000,       // 2
            -0.7070,  0.7070,       // 3
            -1.0000,  0.0000,       // 4
            -0.7070, -0.7070,       // 5
             0.0000, -1.0000,       // 6
             0.7070, -0.7070        // 7
        };

        default : super.plane = {
             0.7070,  0.7070,       // 0
            -0.7070, -0.7070        // 1
        };
    endcase
endfunction

