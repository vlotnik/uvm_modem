//--------------------------------------------------------------------------------------------------------------------------------
// name : pkg_sv_demodulators_types
//--------------------------------------------------------------------------------------------------------------------------------
package pkg_sv_demodulators_types;
    typedef struct{
        int i;
        int q;
    } t_iq;

endpackage