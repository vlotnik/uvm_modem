//--------------------------------------------------------------------------------------------------------------------------------
// name : sincos_envr_cfg
//--------------------------------------------------------------------------------------------------------------------------------
class sincos_envr_cfg extends uvm_object;
    `uvm_object_utils(sincos_envr_cfg)
    `uvm_object_new

    virtual sincos_bfm              sincos_bfm_h;
endclass