//--------------------------------------------------------------------------------------------------------------------------------
// name : tb_complex_multiplier
//--------------------------------------------------------------------------------------------------------------------------------
`timescale 100ps/100ps

module tb_complex_multiplier;
//--------------------------------------------------------------------------------------------------------------------------------
// settings
//--------------------------------------------------------------------------------------------------------------------------------
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // main test package
    import pkg_compmult::*;

    // main settings
    parameter                           A_DW = 12;
    parameter                           B_DW = 12;
    parameter                           TYPE = 0;
    parameter                           PIPE_CE = 0;
    parameter                           CONJ_MULT = 0;

//--------------------------------------------------------------------------------------------------------------------------------
// clock generator
//--------------------------------------------------------------------------------------------------------------------------------
    bit clk = 0;
    // 100 MHz
    always #5 clk = ~clk;

//--------------------------------------------------------------------------------------------------------------------------------
// interfaces
//--------------------------------------------------------------------------------------------------------------------------------
    compmult_bfm #(
          .A_DW(A_DW)
        , .B_DW(B_DW)
    )                                   compmult_bfm_h();

    assign compmult_bfm_h.iclk          = clk;

//--------------------------------------------------------------------------------------------------------------------------------
// DUT connection
//--------------------------------------------------------------------------------------------------------------------------------
    complex_multiplier_wrap #(
          .g_a_dw                       (A_DW)
        , .g_b_dw                       (B_DW)
        , .g_type                       (TYPE)
        , .g_conj_mult                  (CONJ_MULT)
    )
    dut (
          .iCLK                         (compmult_bfm_h.iclk)
        , .iV                           (compmult_bfm_h.iv)
        , .iA_I                         (compmult_bfm_h.ia_i)
        , .iA_Q                         (compmult_bfm_h.ia_q)
        , .iB_I                         (compmult_bfm_h.ib_i)
        , .iB_Q                         (compmult_bfm_h.ib_q)
        , .oV                           (compmult_bfm_h.ov)
        , .oC_I                         (compmult_bfm_h.oc_i)
        , .oC_Q                         (compmult_bfm_h.oc_q)
    );

//--------------------------------------------------------------------------------------------------------------------------------
// UVM test
//--------------------------------------------------------------------------------------------------------------------------------
    typedef compmult_test_default #(
          A_DW
        , B_DW
        , CONJ_MULT
    )                                   compmult_test_default_h;

    initial begin
        uvm_config_db #(virtual compmult_bfm #(A_DW, B_DW))::set(null, "*", "compmult_bfm_h", compmult_bfm_h);
        run_test();
    end

endmodule