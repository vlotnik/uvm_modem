package pkg_logo;
    int nof_logo = 1;

//--------------------------------------------------------------------------------------------------------------------------------
// print logo
//--------------------------------------------------------------------------------------------------------------------------------
    function void print_logo(int logo_sel);
        if (logo_sel == 0) begin
            $display("\t");
            $display("\t                                                                             ...                                 ");
            $display("\t                                                                          .##..##..                              ");
            $display("\t                                                         ....     .......##......###..                           ");
            $display("\t                                                       .###.   ..##....###...........###..                       ");
            $display("\t                                                      .#.###..##........................##.                      ");
            $display("\t                                                     .#..................................#..                     ");
            $display("\t                                                     .#..........####....######...........##..                   ");
            $display("\t                                                     .##.......##.....###.....##............##.                  ");
            $display("\t                                                    .####....##.................##..#####....##.                 ");
            $display("\t                                                    .#...##..............................##...##.                ");
            $display("\t                                                    .#..#...................##...........##....##.               ");
            $display("\t                                                     .##......................#..........##....##                ");
            $display("\t                                                    .##...............................##.......##.               ");
            $display("\t            .######.                                ##....###......#..................#.##....##.                ");
            $display("\t          .#.......#.                              .#.....##.....##......#####.........##.#...##.                ");
            $display("\t         .#.......##                              .##...........##..........##........##.#.#.##..                ");
            $display("\t        .#........#.                              .#..........##.....................##.#.#####.                 ");
            $display("\t        .#.......#.                               .#..........##.......................#.#.###.                  ");
            $display("\t        .#.......#                                ##...........##.....................#...###.                   ");
            $display("\t         .#......#.                               .#....#...............#................###.                    ");
            $display("\t     .....##......#..                             .##.##.###.........######...............##.                    ");
            $display("\t .###....#####......#..                           .##..#.#..  .....   ...###..............##.                    ");
            $display("\t.#.............##....##.                          .###.....####....####...#..............##..                    ");
            $display("\t.#...............##...##..                         .##..............................#####..                      ");
            $display("\t .#..............##....#####..                      .##.......###.................###.                           ");
            $display("\t .#.......####...##....##########...                 .###.......................###.....                         ");
            $display("\t.#.............##......####.....###########################...................######..                           ");
            $display("\t.#...............##...##.##.............................#####..............##..#.....###..                       ");
            $display("\t .#########.......#..##..##............................##....###.............##......##.###.                     ");
            $display("\t .#.........######....#..####..........................##.....######.....####.......##.....###.                  ");
            $display("\t .#.............##...#...######.........................##.......########..........##........###.                ");
            $display("\t  ###..........###..#...############.....................##......................###...........###..             ");
            $display("\t   .############..##..######################..##.........###..................####...............###..           ");
            $display("\t     ..##########...############################.........##..............######....................###..         ");
            $display("\t           ....#############################.##.........##..........#####............................###.        ");
            $display("\t                     ................       .##.........##..........##.................................##.       ");
            $display("\t                                            .##........##..........##...................................###.     ");
            $display("\t                                            ##.........##..........##.....................................##.    ");
            $display("\t                                           .##.........##..........##......................................##.   ");
            $display("\t                                           .##........##..........##..............####......................##.  ");
            $display("\t                                           .##........##..........##.............########....................##. ");
            $display("\t");
        end
    endfunction
endpackage