//--------------------------------------------------------------------------------------------------------------------------------
// name : sincos_agnt_cfg
//--------------------------------------------------------------------------------------------------------------------------------
class sincos_agnt_cfg extends uvm_object;
    `uvm_object_utils(sincos_agnt_cfg)
    `uvm_object_new

    virtual sincos_bfm              sincos_bfm_h;
endclass