//--------------------------------------------------------------------------------------------------------------------------------
// name : raxi_bfm
//--------------------------------------------------------------------------------------------------------------------------------
interface raxi_bfm #(
      DATA_WIDTH = 10
);
//--------------------------------------------------------------------------------------------------------------------------------
    bit                             clk;
    bit                             valid;
    bit[DATA_WIDTH-1:0]             data;
endinterface