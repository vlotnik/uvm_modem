package pkg_demo_basemod;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "common_macros.svh"

    import pkg_modem::*;

    import pkg_vrf_dsp_bfm::*;
    import pkg_vrf_dsp_components::*;
    import pkg_vrf_dsp_modulators::*;

    `include "demo_basemod_test.svh"
endpackage