//--------------------------------------------------------------------------------------------------------------------------------
// name : sincos_bfm
//--------------------------------------------------------------------------------------------------------------------------------
interface sincos_bfm ();
    bit                             iclk;
    bit                             iv;
    bit[11:0]                       iphase;
    bit                             ov;
    bit[15:0]                       osin;
    bit[15:0]                       ocos;
endinterface