`timescale 100ps/100ps

module tb_test_zero_project_top;
//--------------------------------------------------------------------------------------------------------------------------------
// libraries
//--------------------------------------------------------------------------------------------------------------------------------
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "common_macros.svh"

    import pkg_modem::*;
    import pkg_demo_basemod::*;

    `print_logo

//--------------------------------------------------------------------------------------------------------------------------------
// clock generator
//--------------------------------------------------------------------------------------------------------------------------------
    bit clk = 0;
    // 100 MHz
    always #50 clk = ~clk;

//--------------------------------------------------------------------------------------------------------------------------------
// interface
//--------------------------------------------------------------------------------------------------------------------------------
    if_ddc_bfm #(.INCH_NUMBER(2)) if_ddc_bfm_h();

    assign if_ddc_bfm_h.clk         = clk;
    assign if_ddc_bfm_h.iq_v        = 1;

//--------------------------------------------------------------------------------------------------------------------------------
// UVM test
//--------------------------------------------------------------------------------------------------------------------------------
    initial begin
        uvm_config_db #(virtual if_ddc_bfm #(.INCH_NUMBER(2)))::set(null, "*", "if_ddc_bfm_h", if_ddc_bfm_h);
        run_test("demo_basemod_test");
    end

//--------------------------------------------------------------------------------------------------------------------------------
// dump
//--------------------------------------------------------------------------------------------------------------------------------
    bit dump_v;
    bit[15:0] dump_i;
    bit[15:0] dump_q;

    assign dump_v = 1'b1;
    assign dump_i = if_ddc_bfm_h.iq_i[0];
    assign dump_q = if_ddc_bfm_h.iq_q[0];

    `dsp_dump_to_file(4, dump, dump_v, {dump_q, dump_i}, clk)
endmodule