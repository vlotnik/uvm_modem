//--------------------------------------------------------------------------------------------------------------------------------
// name : pkg_modem_math
//--------------------------------------------------------------------------------------------------------------------------------
package pkg_modem_math;
    real c_pi = 3.1415926535897932384626433832795;

    function real f_abs_real(real x);
        real result;
        result = x < 0 ? -1.0 * x : x;
        return result;
    endfunction
endpackage