//--------------------------------------------------------------------------------------------------------------------------------
// name : raxi_bfm
//--------------------------------------------------------------------------------------------------------------------------------
interface raxi_bfm #(
      DW = 10
);
//--------------------------------------------------------------------------------------------------------------------------------
    bit                                 clk;
    bit                                 rst;
    bit                                 valid;
    bit                                 ready;
    bit[DW-1:0]                         data;
endinterface