package pkg_demo_basemod;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "common_macros.svh"

    import pkg_vrf_dsp_components::*;

    `include "demo_basemod_test.svh"
endpackage