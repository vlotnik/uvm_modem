//--------------------------------------------------------------------------------------------------------------------------------
// name : pkg_rounder
//--------------------------------------------------------------------------------------------------------------------------------
package pkg_rounder;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "common_macros.svh"

    import pkg_modem_math::*;

    import pkg_raxi::*;
    import pkg_pipe::*;

    `include "sim_rounder.svh"
    `include "rounder_scrb.svh"

    `include "rounder_base_test.svh"
endpackage