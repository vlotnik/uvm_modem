//--------------------------------------------------------------------------------------------------------------------------------
// name : tb_sin_cos_table
//--------------------------------------------------------------------------------------------------------------------------------
`timescale 100ps/100ps

module tb_sin_cos_table;
//--------------------------------------------------------------------------------------------------------------------------------
// settings
//--------------------------------------------------------------------------------------------------------------------------------
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // main test package
    import pkg_sincos::*;

    // main settings
    parameter                       FULL_TABLE = 0;
    parameter                       PHASE_W = 12;
    parameter                       SINCOS_W = 16;
    parameter                       PIPE_CE = 0;

//--------------------------------------------------------------------------------------------------------------------------------
// clock generator
//--------------------------------------------------------------------------------------------------------------------------------
    bit clk = 0;
    // 100 MHz
    always #5 clk = ~clk;

//--------------------------------------------------------------------------------------------------------------------------------
// interfaces
//--------------------------------------------------------------------------------------------------------------------------------
    sincos_bfm                      sincos_bfm_h();

    assign sincos_bfm_h.iclk = clk;

//--------------------------------------------------------------------------------------------------------------------------------
// DUT connection
//--------------------------------------------------------------------------------------------------------------------------------
    sin_cos_table #(
          .g_full_table             (FULL_TABLE)
        , .g_phase_w                (PHASE_W)
        , .g_sincos_w               (SINCOS_W)
        , .g_pipe_ce                (PIPE_CE)
    )
    dut(
          .iCLK                     (sincos_bfm_h.iclk)
        , .iV                       (sincos_bfm_h.iv)
        , .iPHASE                   (sincos_bfm_h.iphase)
        , .oV                       (sincos_bfm_h.ov)
        , .oSIN                     (sincos_bfm_h.osin)
        , .oCOS                     (sincos_bfm_h.ocos)
    );

//--------------------------------------------------------------------------------------------------------------------------------
// UVM test
//--------------------------------------------------------------------------------------------------------------------------------
    initial begin
        uvm_config_db #(virtual sincos_bfm)::set(null, "*", "sincos_bfm_h", sincos_bfm_h);
        run_test();
    end

endmodule